module top_module( input in, output out );

    // This is a NOT gate
    // ~ is the not/invert operator
    assign out = ~in;

endmodule
