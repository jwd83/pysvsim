module rom_deadbeef (
    input  logic [1:0] addr,
    output logic [7:0] data
);
    // ROM data loaded from deadbeef.txt by simulator
endmodule
